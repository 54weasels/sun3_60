$ 3bitcom
$ JED2CKT -- JEDEC File to OPALsim Circuit/Macro Translator (Version V055)
$ Copyright (c) National Semiconductor Corporation 1990,1991
$ Translated from 3bitcom.jed. Date: 3-20-92
$ DEVICE GAL16V8
$ PERIOD 20

.LIB 3bitcom.mac

* U1 3bitcom 2 a2 a1 a0 nc compare nc b2 b1 b0 GND nc nc lt nc
+ eq nc gt nc nc VCC

a2 INPUT 0 20 = LLHHLLLLLLLLLLLLLLLLLLLLLLLLLLLL
a2 INPUT 760 20 = H
a1 INPUT 0 20 = LLHHHHLLLLLLLLLLLLLLLLHHHHHHHHHH
a1 INPUT 760 20 = LLLLLLLLLLLLLLLLHHHHHHHHHHHHHHHH
a0 INPUT 0 20 = LLHHHHLLLLLLLLHHHHHHHHLLLLLLLLHH
a0 INPUT 760 20 = LLLLLLLLHHHHHHHHLLLLLLLLHHHHHHHH
compare INPUT 0 20 = HLHLHLHHHHHHHHHHHHHHHHHHHHHHHHHH
b2 INPUT 0 20 = LLHHHHLLLLHHHHLLLLHHHHLLLLHHHHLL
b2 INPUT 680 20 = HHHHLLLLHHHHLLLLHHHHLLLLHHHHLLLL
b2 INPUT 1320 20 = HHHH
b1 INPUT 0 20 = LLHHLLLLHHLLHHLLHHLLHHLLHHLLHHLL
b1 INPUT 640 20 = HHLLHHLLHHLLHHLLHHLLHHLLHHLLHHLL
b1 INPUT 1280 20 = HHLLHH
b0 INPUT 0 20 = LLLLLLLHLHLHLHLHLHLHLHLHLHLHLHLH
b0 INPUT 640 20 = LHLHLHLHLHLHLHLHLHLHLHLHLHLHLHLH
b0 INPUT 1280 20 = LHLHLH

.BUS seta a2 a1 a0
.BUS setb b2 b1 b0

.PROBE compare seta setb lt eq gt

.TIME 1399

.END
